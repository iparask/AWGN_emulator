library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity myrom2 is
port( 
	  address1	: in signed (9 downto 0);
	  address2	: in signed (9 downto 0);
	  address3	: in signed (9 downto 0);
	  address4	: in signed (9 downto 0);
	  stoixeio1	: out signed (31 downto 0);
	  stoixeio2	: out signed (31 downto 0);
	  stoixeio3	: out signed (31 downto 0);
	  stoixeio4	: out signed (31 downto 0)
);
end myrom2;


architecture struct of myrom2 is

    type rom_type is array (623 downto 0) of signed (31 downto 0);
    constant stoixeia : rom_type :=( "00111010111111000001000111000110","01010111111001101011001001000110","11101001111101010110110110101110","11001100011100001101011100000001","00001101111100110100001001010011",
"11101001000011010001000010100001","10001101101110011100001011111101","11110010110111100000011101110010","01001100110101011111000100010101",
"10111000001000001011101101010100","01100010110000011110011010100000","00101001001010011111111101100001","01110011011000100100011001000100",
"01101111111000001100011111010001","11001001011010101000001110111110","10001000101001100101010100100000","11111110001101101111111011100001",
"01000001010001011110111100110011","00110100000000000101101101101010","10100100011010011101011010101101","11010010111010100001110110110110",
"10010010010101101011100100001001","10100110110000111001111100100100","10010011100100000010101000000000","10000101111000000011011001101101",
"11100111111101101001001101010111","01111100001100011101111011010010","01100110101100110101011100011101","11010100101100100111011001101110",
"11111011100011111101110001110000","01000111001000010001000011100001","10110000010001011010000000010101","01110010011001111100111100000100",
"10001001010110011100110111001011","11001011010110110001101110010001","11101000011110011010010110101111","10011100111010100010110100010101",
"00101001001010001010000010101110","11000110010001111011010100000010","10111101110000001000011110000001","11101011111101000111001110100011",
"00001100001111010000101100110000","01100101011001110100110101110101","00111011000001010010011101101000","10110111011100001100011100100110",
"11001100111110001001001101010001","01010100001010101011000001100101","01000001101111110000101100001011","10001010000010101110100000011110",
"11011000100010100000111010101001","11010110111000001010100101110111","11100001111110101100001010110111","01001011111100011000011111010110",
"01100110100110001001111000111001","10111100001111100000101010000100","10010001010010101000011110011000","10100101011110110000000010000101",
"10010010111110111000110001011101","01001100100010101001101101000101","11110001101011001001000110000011","01111001101010001011111000001100",
"11101011101110101101111000100001","11101111000101101011101010001111","01101111000111111001001101111101","10000101001110001101011101000111",
"11000101000111010000000001011101","00110101000100000001000100111100","10101010011000110101010101001001","00000101010111101100011001111100",
"11010100010111001000111011100010","01110011100100001000001011101010","01100010000111100001100100110111","10001101101101000110010110111100",
"10011110011001011101100001110110","01101010100011101011101110110000","11001100100001101110001011100001","01000001001101001111000000000111",
"10000010100011011011001001000100","10111000101001110100101000010011","00000101101111010001110101001111","10010101100001011001011100101110",
"01101100001100001010011001101100","00000000010010100111010000100001","00101000000011100010100011000101","00111001111100011010001011010010",
"10011000010110101010011111000110","01001010011100111000110000010010","11110011100110111010000010101100","01010001100000011111001001100111",
"10010001000110000000101110001011","00101110001010011001011011011001","00010000111101011011001010000110","01001110101011101110110000001010",
"10011001010101011100100101010100","10100010111011111111011101101001","01110001110001001100001111000110","00110101100101111111001000001000",
"11100011101010000100111011010000","11111010001010110110000010011101","00101001011011001101011100100111","01010000111101100001110001101100",
"10001100010110101000101110010110","11111111010001011000010110010000","11110101100011000101111110110111","10001011010101011101100100001100",
"01111010011000110100011110111000","01110011101010010111111011001111","11001011010011110011101101101111","10110100101000110110110100100001",
"10011101000001111001111011110100","11000010010111101010101001110011","01001010111010010110101000111000","11111000010100110000001000000000",
"10110100111001110010101001010111","10000001001111111010100101110101","10110101101001100100111000110011","10010010000000010110111000101101",
"10101001001000001011011010101100","10101110101110001011001100111100","01001101110000011010010000000100","10110101111111101101001011101000",
"01000110110111101101010101111110","01000111001011000011101001110111","10011011000000000000100110101000","11101011001001001111110111110000",
"11011011000100111010101111001000","01110111100010011001101001110011","10110010100110010010101010110001","01010100000010011101000000011101",
"11100101010001010011111001010101","11011001111111011110010010111101","01010100000011011001101111010100","01001110010011010100100100111000",
"00000010010100011011000001110010","01011100000000000011101010100111","01011101001111011110111101101000","11111011100101011000010000001111",
"10011110010110110011110011101011","01100010010101011111001010010001","10101011010010001101110011111010","00010111111001111100010001110100",
"01101101000001001000001011100000","00011000101110000100110110100000","11001100001100101101001100000111","01100111001011101011111011011001",
"01100101110010110100100001010001","01110101001001111010111100011000","00011011110000011011000010000101","11111100010100110111111001100110",
"11110000000110101110101100000001","01100100011110000000110011011011","10101111100111000001001111111110","01101101011010110010100001000110",
"01110100000001110010101101010010","10000101011000110011100110010110","11000000011011110011011001100000","01111011011111100011000110101000",
"10011011011110011100001110010110","00011010110001100100100011100111","11101001010101011011001000100101","10100000110010011000011001111000",
"11101000010111000111001111101010","01110110100101111010011101110100","10110011011110110001110101001100","00001001100001011100111010010000",
"10100010010101000011001100000011","01110000110101010111011101000001","01011001110000100001100110101110","00110100100110101111100100101110",
"11000001101000001000111001101101","00100000010000110010100100010111","00001111110101110100000001100011","01001110100111100110110000010001",
"10011111110011101001101100000001","00010101001101010101001000100010","01001010011111001100010010101100","10111001101011111111011100110000",
"01111100011110010100110010011001","01101111010101110010100001001011","01100111111101111111010101000001","01000011110101010000100100000001",
"11000011110000101100000000000101","11101010111011001011110010011110","00111000000000011000111011101111","11001010001110011101111000011110",
"00110110000111110111111100010110","00011001010111110011010101111111","00110111111100100010001101010111","01000101000101101001000010101100",
"10100101111000111100110100111010","10100110100100100110011111010010","00011001111110101010111001000101","10001100110010110001010011110111",
"01000111100100111111000000100100","01110110111101001100111011101001","10101110010000001011101001010100","11001000110101101111010111011000",
"00110101010000001110011011001110","01101001111100011110110011111011","00001100110111101100101001001010","11010110111010010111110100111001",
"01100001100100111001001001011111","01101110101001001110000100000111","10101110011011011100001111011010","01000101101111001000000101011111",
"01011001001000011000110110011011","11101111100110101000011001110111","00110011110110000000001001111000","00000111101010000100000011111111",
"11001001111111001111101110011100","00111100101001101100111011100110","11101010000101111011000000001011","10111100100000101011101110101111",
"10001001001010001111010111001000","11000001100110011111000010001010","00101100101111001100101111001000","10000011111111111101101101000110",
"01110001101001001001110101011001","00110111100111111111111001010101","10010111100111110100111111111011","00010011111110011111100100010111",
"11010001000001001101011111111101","10000011110010000110000100110100","00101111000010111110000110100011","10000111000100000100101010101111",
"11101111011000001111111011001001","11010000001010101111100110011111","00001000011010101000100011001110","01010010011000111100101110111010",
"10011111100100010011001111110101","11110001111010010101010100111000","10010010011101010110000100011010","00111010111000011110100111100000",
"11101101101110000011011001000110","00000010111111011001000001101101","11001001100001110111101011100000","00111101010000001111110010100110",
"01000000110111011010011111011101","10101101011001011110101011010110","01001011001010001111110110101010","11101000110001000001100111101010",
"11010011011101111111110001110000","00111110110001010110010010010010","10101011011001000110111010100011","00010011111100010010101110001111",
"00111110111111101110001001011010","10001000011001100101010101111011","00000010110011001001100110100101","01100110101100110100010010001111",
"10110010010100111011111101000011","00010001011001100010101010011010","11001010101001011000110010110101","00000101111101010111011000111110",
"00011000000011001110001001111100","10110111000111010001100011010001","01010110110010111011011000010001","01000100011010111101011001111100",
"01010111011101011000001111110011","01100011001001101111100111011101","00110011100000110111000110101100","11100011001010101100010101011011",
"11011111100111110100000111100001","01011011110110111011011110011010","10000010010011101001001110011001","00100100001111010100110111000001",
"01111110110100110010110000101000","01100011011010001011010101111001","10000011101101110100010001100011","11001110110000101100010010110001",
"11100100100011000110010111110001","00001001010000111101011101011010","00110001000011010100101010010110","11000001100101111001010100101001",
"00110010000101010110011101101000","00111011001101011011010101011111","11101010110011111011000010101101","00100000001101110100101110101111",
"00111100001011110011101010011000","11111001001101001000100100011100","00110000111110101000011011000111","11000000011100011100110111101110",
"10011111011000010011100100001001","11000101000101111110101100100100","01000100011000001010100010100100","01010000100111111011111010111110",
"00010100100100111001110011101110","01000001100000000111001100101110","00000111110100001011000000100110","10110100000111011111010000000100",
"10111111100100101000100111111001","01000011101101010011111101101101","11000001111000000100101000011001","11000000100000010001001100100001",
"11100011101111111010100000010101","11111110110111101011011010100110","01100001111100010001011110101011","10011111010100100111100001111101",
"11011101010000001111010011011100","00001011100111111101110010110010","11010000011110001110010111110100","00001000111000000101111000000010",
"00000110010100001101010100001101","11110010001101000001101110011011","11110100111010111011011000100010","11010111001000000010001011010000",
"10000101100110100100111011100011","11101101010001101001011001101100","10101000001011101000011011011111","10010000110010000111001101000001",
"11100101010101111000110111101111","10000010100101100011111110011101","10101100100010110101000001011000","00000111100000001011111000101001",
"00011101000100001101100001000011","01100011110011011001111110111110","01010101100011010101010011011000","01110000010001010011000001001100",
"01001110111011001000100011000000","01100011010101111000101001110010","01001000111000100011101111010011","00000010000100100111001101100011",
"11101010010011001111101110100100","01110010010000000101110001011110","11111111010011011100101110010010","10100000010010000001111001110001",
"00001110011010011001110000000010","00101000000100100000000100100001","11001111011001000110001010100101","11000001001110000110000011001100",
"01100110100100010111010000000110","01110101001001011100110010000111","01001110011100100000001111101111","10010100101000010101111110011011",
"00010100001011001000011011001010","00001001100110011100011001110110","00101110010101000011001110110010","10011100111011110011100110110010",
"10011011100111101111010010011001","01110001011110101101010010011100","01111001001011111000110010111000","01111111000111010111010001111011",
"00011010101011011101111011101010","11101000111100000011010100100010","11100100100111001111010000010011","01010010000000011011000110011100",
"01000011010110100010110110100001","00001011100000110000111000001110","00110101010111100100001101100011","11100101010100110000010000011110",
"11010000010010111010011010010101","00001111010110101010110000111001","01001000001111010101111110111010","01011110110100111010110110001011",
"10000011000001100011011100111100","11010111101001101001011101100100","01001010110111010110010010000101","11101110100111101011110111110010",
"11101010111101001111100101010001","11100100010110101011000001111110","11011110101111001100000111101000","00110011001100001011011110111011",
"11101101000011100111100000011011","01111100101011000001111001011000","10111010011011010101100100101101","10110001101001110100110010111101",
"11001000110011010110110100011000","00010011001100001100111011100000","11001100001100011010100110101001","01011001001111111001010011001111",
"00101000000010111001111111110001","11010011100100100110101011111110","11011110001111111000001011011100","11001011000010111110011010001101",
"11010100101001110111111001011110","00111011111001011010010011101000","00001101110010101110111101100100","11000100111101101010000101111011",
"01101100001001100001011111111110","11010000100000000111110110010100","00111010111011110010101000010011","00111101110001110011011110000100",
"01100110100111011100010000111101","00010000010000101011000101111111","10111011001001010011110011000001","11100101011000111110111100111011",
"10011010011011010101001110001110","10000010111111010001001111011011","01100010000100011011110100001100","10010110110111011110111001010110",
"01110100011001001110000011110111","11001111000010101100101011000010","11100011101011011100100000001010","01000101110000110011000000110000",
"11111010100001001000111100000100","10101110110100001111001001111101","01010110110101100010110000001110","10110000100111010111101011100000",
"10111100001110101010101010111110","10011011010110011001100100111110","10001111001111110000010010000010","00110110000101101011000001011011",
"11001110001000111011111100001110","00101000001011110011110111100111","00101100101100000011000111001001","11010101000111011011001101011110",
"01100100111000100001010010100000","01010101101001110101111100100001","00010000000010000000110110110110","11001001101011001011001111110011",
"01011110001111010100110101110011","01001111010001100011110100101001","10000001111111110010100011000001","00110000101011000010110101001111",
"00011100111100011010011000010010","10101111000001111001001100111010","10110110110101000010000100001110","01110001000110101001101000100100",
"01001110101010010010001110010010","00001011110001011001110010010110","01010011001111010111011101000111","01011011000010100101000001100000",
"11111011110010101011011111110010","00011100010000010010011000100010","11110010111111110001000000101100","01110110101100010000111000100011",
"10101111100111010101101100100110","11001000101001111000001111111111","10100111011111101101110010101011","11101110101011100000000001011111",
"10011111000111101000111110110000","00100000110000001111101010110010","01011011100110111010001100000011","11010001101101101000111111101111",
"11100100101100111101100111000011","10110110111011100100101010110111","00010101000010110001010100001101","00011101011000010010010010001011",
"01011011000011000111001011110010","11110110011111011001001010110100","11110001011001111110011001011110","01100101000100101110100000010010",
"10011010101001101100010000011010","00010110010011010011001111110101","10001110000000110111101011111100","01000101111111010110001001011110",
"01111110110001111110111011111001","10011011000100010110111011000000","10000001011111001110011011001000","10100011101000010100100110110001",
"01101111101100110011111111011111","10000110111101000111101000110101","01100001111011011011111011000111","10011000010100001001001010110010",
"00110111010000110110111100100101","10101010101110010000110100000101","11000000000111001110101011111011","10011110100011100010000011001011",
"01110001101001110001100110110000","11000000000111101011011001010110","01111110011100011100010100111100","01001100111000110001111111100111",
"01110110100110111110011111110001","00101111100011000111001101001100","01011010101111000110111011101011","00110011101101111011000100111000",
"10100101100110000101101011000001","00110000110011101010110101111100","01011010011110110001101110011110","10110010111110010000100101111101",
"11010101010110011011111110101001","11001100111101011110010010101000","00100010100100111010000100100101","00010110000010110001111010001010",
"10111010100111000011111111101100","00000001111101001100110001100011","01011000110011000010100100100011","00101110100101100100011010001001",
"01111000000011010010111000001111","01101101111000111100001011001110","10110101101100111110010000010001","01011100101111110111110001010100",
"11001111000010010000101100011110","10101010010101010000100000000101","10110100101111011010101101100000","11010010001010001001110010100000",
"01001000000101011110000101001110","11001110110000111001000101101000","00011001010011111010100110111111","01101111011111101100000111110011",
"10101110001001100101100111000101","01101011101000110001001101000011","10011100100110100111110011100110","00111100101011011010011100000111",
"11010011010011010010010110010000","00011100111100101000111001101111","10110111111100110000110111100110","10011110111100111100111011010011",
"10001111011101010001101010011000","00111100111000101111111100011000","10100111101011101001100010000001","11100000100101100110111010000001",
"11001100111011010100111010000101","11110010001001001011110100110101","11010111000101001001010000100110","00001011011001001100000000111010",
"11101101011001101001110101101000","00101100010000101110100110010101","00111011100000010001011100011100","10110011101011111010111000011111",
"01110101101101011100010101100101","10011100100001100001111001111110","00100111000011110011110101010101","01101101111111101011010010010000",
"00000011110001110100110101010011","01000000011101011111000100011001","01010110000011001011000110011001","10001111001110001010101000110111",
"01010100111010110010110101011100","11100000101110101001101000110111","01001000000000001101101111010101","11110101001001100011010011100001",
"01000011011100110010011101111101","10111000100010001000101100011001","00110111101110101110001111111010","00011001100010011110111011110000",
"10110011001110000111101101111110","11011101010011001111110101111110","11011001000110011000001111110100","10101111011110110011011011010101",
"00000101111101000011110001011111","10000110111101000110001101011010","01110111010010000100111101010111","01100010100010101011000101000101",
"11001011010101100000110010111110","11001011110110101100000000011001","11111010011001110100001010111001","10010100001010010101101111110010",
"11111111110000001011111000011011","00111100000011010010011011011100","10010110000110011000110011000000","10001100101011100001101010010110",
"11111101010101010110000010111110","11101001010011011001010001110101","10110011011011001100110100010001","01010010110111111011010001011001",
"00110101111111111110101101111000","01011010100010111010101110000011","01001011011101011111100110100101","01011010000011111110001011101111",
"10001011111111000000011101011100","00100010110001011101010101011110","11000000000110101111111000010101","10010001000001101110100010000001",
"11001001001011011111011101111001","11100011101111010110011111111010","00000001111110101111010011101110","00110001111001111110011000100010",
"10011010000101001111011000101001","01000111110100011101011110011011","01100011111010101000001010100111","00110110001001010001101100100011",
"10000100101011110010110010100010","01000000010101111111011111000010","01011111010111001000001110111101","10011111010001011011011100111000",
"00010010001111110110000101101011","00010111001000011101001000001110","01001111000110101001001100100111","01001011110001111110000100101011",
"10110110100110000101100100001001","01001011000110100110111010010011","11100100111010111100001111100101","11110110100100110111001110100111",
"11101000011110101101100001100100","00100001110101101100101101101101","10101110011010000011010110001110","01111010011101110010010010001000",
"01101100100110010110001010010001","00010101101010001001000010010100","10010101101000111101111011001111","10000011001001000010100100110010",
"11111001110010010011101011101011","00100011110001001010101111101001","00101111100011111001001101111101","11101011011110001000100010010100",
"00100110001011100000101110011110","00010101111110100001010010001110","10011111110010101001101101011110","11011011100110010010010000100101",
"00100010000110100001011010001101","10001110110000010111010100101101","01010101111111001100000110000000","00110111101111110100100100110101",
"10101100011000001001101100111001","11101011111010101011100100111101","00101000011001001011111010011000","01001111000101111100110011001111",
"01000101000110010101010011001010","01011000010010111011101001100001","00000110101001001000001000101000","10000000110111101101011101001010",
"01011000010100001011001011010101","00000010110001001111011011111011","11000100001111111010100001101100","11100001001011011111000011000101",
"10100010010110000101010000000100","01001111010111100110011111001011","01010000010000100111100101110101","00110000001110111100011101010010",
"10100100101100101011000101100001","00001010100111010111001101111000","10010010110111000011101101101010","10010000010110111100111111111110",
"10001001001110010111011000101000","00111010111010010100010110000111","11001011001010110110111110000110","10101100000101010111000110000110",
"10010111010100110110010000001001","00011011111000000000010001010110","01110111101010000001001010011001","11001001110000010111010011100010",
"00100000011100000110111011010101","10000111111001111000100110101100","11010111100110000011111011001110");  

begin

stoixeio1<=stoixeia(to_integer((unsigned(address1))));
stoixeio2<=stoixeia(to_integer((unsigned(address2))));
stoixeio3<=stoixeia(to_integer((unsigned(address3))));
stoixeio4<=stoixeia(to_integer((unsigned(address4))));
end struct;
